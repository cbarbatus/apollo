@media screen and (min-width: 671px) {

    body {background: url(/img/rcg_large_text.png) no-repeat,
            url(/img/newtree1920.jpg) top center no-repeat;
        color:black;
        font-family: font-family: 'Cabin', sans-serif;
        font-style: normal;
    }

    .startpad {
        position: relative;
        top: 160px;
        width: 100%;
    }
}



body {
    background-color: #296523;
    font-family: 'Cabin', sans-serif;
    color: black;
}

.embed-container {
    position: relative;
    padding-bottom: 50.625%;
    padding-top: 30px;
    height: 0;
    overflow: hidden;
    max-width: 90%;
    display: block;
    margin-left: auto;
    margin-right: auto;
}

.embed-container iframe,

.embed-container object,

.embed-container embed {
    position: absolute;
    top: 0;
    left: 0;
    width: 100%;
    height: 100%;
}

.btn-go {
    background-color: #67b168;
    border-radius: 8px;
    font-weight:bold;
    color: #000;
}

.btn-warning {
    background-color: yellow;
    border-radius: 8px;
    font-weight:bold;
    color: #000;
}

.btn-danger {
    background-color: red;
    border-radius: 8px;
    font-weight:bold;
    color: #000;
}

.btn-go:hover,
.btn-go:focus,
.btn-go.focus,
.btn-go:active,
.btn-go.active,
.open > .dropdown-toggle.btn-info {
    color: #ffffff;
    background-color: #4b914b;
    border-color: white;
    text-decoration: none;
}

hr {
    border-top: 2px solid #000;
}

table {
    background-color: #e0f2ff;
}

td, th {
    padding-left: 4px;
}

blockquote {
    background-color: #f8f8ff;
}

li {
    font-size: 100%;
}

a {
    color: #0000ff;
}

a:hover, a:focus {
    color: #8888ff;
    font-weight: bold;
}

.tab { margin-left: 40px; }

.TextWrapRight {
    float: right;
    margin: 10px;
    clear:left;
}

.TextWrapLeft {
     float: left;
     margin: 10px;
     clear:right;
 }

img.bordered {
    border:groove black 4px;
}

.navbar {
    padding: 0rem 1rem;
}

.card {
    background-color: #dcf0ec;
}




.note {
    font-style: italic;
    color: darkred;
}

h3, h2 {
    font-weight: bold;
}

.dropdown-item:hover,
.dropdown-item:focus {
    color: white;
    background-color: #343a40;
}

.dropdown-menu {
    color: white;
    background-color: #343a40;

}

.dropdown-item {
    color: white;
}

